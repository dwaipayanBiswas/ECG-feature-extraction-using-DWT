`timescale 1ns / 100ps

module ecg_top_stim;

reg [15:0]  data_in;
reg clk, nReset;

wire [15:0] q_peak_ref,q_peak_pos_ref,r_peak_ref,r_peak_pos_ref,
s_peak_ref,s_peak_pos_ref,start_qrs_fin_2,end_qrs_fin_2,
p_begin,p_end,p_peak,p_peak_pos,t_begin,t_end,t_peak,t_peak_pos; 

ecg_top top (q_peak_ref,q_peak_pos_ref,r_peak_ref,r_peak_pos_ref,
s_peak_ref,s_peak_pos_ref,start_qrs_fin_2,end_qrs_fin_2,p_begin,p_end,p_peak,p_peak_pos,t_begin,t_end,t_peak,
t_peak_pos, data_in,clk,nReset); 

always
begin
	     clk = 0;
  #500000	clk = 1;
  #500000	clk = 0;

end

initial
  begin
           nReset= 0; 
		 data_in = 	9;
      #250000 nReset= 1;


#2200000 data_in = 	9;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	17	;
#1000000 data_in =	17	;
#1000000 data_in =	17	;
#1000000 data_in =	17	;
#1000000 data_in =	17	;
#1000000 data_in =	17	;
#1000000 data_in =	26	;
#1000000 data_in =	26	;
#1000000 data_in =	26	;
#1000000 data_in =	26	;
#1000000 data_in =	26	;
#1000000 data_in =	26	;
#1000000 data_in =	26	;
#1000000 data_in =	26	;
#1000000 data_in =	26	;
#1000000 data_in =	26	;
#1000000 data_in =	26	;
#1000000 data_in =	26	;
#1000000 data_in =	26	;
#1000000 data_in =	26	;
#1000000 data_in =	26	;
#1000000 data_in =	26	;
#1000000 data_in =	26	;
#1000000 data_in =	26	;
#1000000 data_in =	26	;
#1000000 data_in =	26	;
#1000000 data_in =	26	;
#1000000 data_in =	26	;
#1000000 data_in =	26	;
#1000000 data_in =	26	;
#1000000 data_in =	26	;
#1000000 data_in =	26	;
#1000000 data_in =	26	;
#1000000 data_in =	26	;
#1000000 data_in =	26	;
#1000000 data_in =	26	;
#1000000 data_in =	26	;
#1000000 data_in =	26	;
#1000000 data_in =	26	;
#1000000 data_in =	34	;
#1000000 data_in =	34	;
#1000000 data_in =	34	;
#1000000 data_in =	34	;
#1000000 data_in =	34	;
#1000000 data_in =	34	;
#1000000 data_in =	34	;
#1000000 data_in =	34	;
#1000000 data_in =	34	;
#1000000 data_in =	34	;
#1000000 data_in =	34	;
#1000000 data_in =	34	;
#1000000 data_in =	34	;
#1000000 data_in =	34	;
#1000000 data_in =	34	;
#1000000 data_in =	43	;
#1000000 data_in =	43	;
#1000000 data_in =	43	;
#1000000 data_in =	43	;
#1000000 data_in =	51	;
#1000000 data_in =	51	;
#1000000 data_in =	51	;
#1000000 data_in =	51	;
#1000000 data_in =	59	;
#1000000 data_in =	59	;
#1000000 data_in =	59	;
#1000000 data_in =	59	;
#1000000 data_in =	68	;
#1000000 data_in =	68	;
#1000000 data_in =	68	;
#1000000 data_in =	68	;
#1000000 data_in =	76	;
#1000000 data_in =	76	;
#1000000 data_in =	76	;
#1000000 data_in =	76	;
#1000000 data_in =	76	;
#1000000 data_in =	76	;
#1000000 data_in =	76	;
#1000000 data_in =	76	;
#1000000 data_in =	76	;
#1000000 data_in =	76	;
#1000000 data_in =	76	;
#1000000 data_in =	76	;
#1000000 data_in =	76	;
#1000000 data_in =	76	;
#1000000 data_in =	76	;
#1000000 data_in =	76	;
#1000000 data_in =	76	;
#1000000 data_in =	85	;
#1000000 data_in =	85	;
#1000000 data_in =	93	;
#1000000 data_in =	93	;
#1000000 data_in =	101	;
#1000000 data_in =	110	;
#1000000 data_in =	118	;
#1000000 data_in =	118	;
#1000000 data_in =	127	;
#1000000 data_in =	135	;
#1000000 data_in =	144	;
#1000000 data_in =	144	;
#1000000 data_in =	152	;
#1000000 data_in =	152	;
#1000000 data_in =	152	;
#1000000 data_in =	152	;
#1000000 data_in =	152	;
#1000000 data_in =	152	;
#1000000 data_in =	144	;
#1000000 data_in =	144	;
#1000000 data_in =	135	;
#1000000 data_in =	135	;
#1000000 data_in =	127	;
#1000000 data_in =	118	;
#1000000 data_in =	110	;
#1000000 data_in =	110	;
#1000000 data_in =	101	;
#1000000 data_in =	93	;
#1000000 data_in =	93	;
#1000000 data_in =	85	;
#1000000 data_in =	85	;
#1000000 data_in =	76	;
#1000000 data_in =	76	;
#1000000 data_in =	76	;
#1000000 data_in =	76	;
#1000000 data_in =	68	;
#1000000 data_in =	68	;
#1000000 data_in =	68	;
#1000000 data_in =	68	;
#1000000 data_in =	68	;
#1000000 data_in =	68	;
#1000000 data_in =	68	;
#1000000 data_in =	68	;
#1000000 data_in =	68	;
#1000000 data_in =	68	;
#1000000 data_in =	68	;
#1000000 data_in =	68	;
#1000000 data_in =	59	;
#1000000 data_in =	59	;
#1000000 data_in =	59	;
#1000000 data_in =	59	;
#1000000 data_in =	59	;
#1000000 data_in =	59	;
#1000000 data_in =	59	;
#1000000 data_in =	59	;
#1000000 data_in =	59	;
#1000000 data_in =	59	;
#1000000 data_in =	59	;
#1000000 data_in =	59	;
#1000000 data_in =	59	;
#1000000 data_in =	59	;
#1000000 data_in =	59	;
#1000000 data_in =	59	;
#1000000 data_in =	59	;
#1000000 data_in =	51	;
#1000000 data_in =	51	;
#1000000 data_in =	51	;
#1000000 data_in =	51	;
#1000000 data_in =	51	;
#1000000 data_in =	43	;
#1000000 data_in =	43	;
#1000000 data_in =	34	;
#1000000 data_in =	34	;
#1000000 data_in =	26	;
#1000000 data_in =	26	;
#1000000 data_in =	17	;
#1000000 data_in =	17	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	0	;
#1000000 data_in =	0	;
#1000000 data_in =	0	;
#1000000 data_in =	-7	;
#1000000 data_in =	-7	;
#1000000 data_in =	-7	;
#1000000 data_in =	-7	;
#1000000 data_in =	0	;
#1000000 data_in =	0	;
#1000000 data_in =	0	;
#1000000 data_in =	0	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	0	;
#1000000 data_in =	0	;
#1000000 data_in =	0	;
#1000000 data_in =	0	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	0	;
#1000000 data_in =	0	;
#1000000 data_in =	0	;
#1000000 data_in =	0	;
#1000000 data_in =	0	;
#1000000 data_in =	0	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	17	;
#1000000 data_in =	17	;
#1000000 data_in =	26	;
#1000000 data_in =	26	;
#1000000 data_in =	34	;
#1000000 data_in =	34	;
#1000000 data_in =	26	;
#1000000 data_in =	17	;
#1000000 data_in =	0	;
#1000000 data_in =	-15	;
#1000000 data_in =	-49	;
#1000000 data_in =	-83	;
#1000000 data_in =	-133	;
#1000000 data_in =	-184	;
#1000000 data_in =	-243	;
#1000000 data_in =	-310	;
#1000000 data_in =	-378	;
#1000000 data_in =	-453	;
#1000000 data_in =	-521	;
#1000000 data_in =	-596	;
#1000000 data_in =	-664	;
#1000000 data_in =	-731	;
#1000000 data_in =	-790	;
#1000000 data_in =	-849	;
#1000000 data_in =	-900	;
#1000000 data_in =	-942	;
#1000000 data_in =	-984	;
#1000000 data_in =	-1018	;
#1000000 data_in =	-1043	;
#1000000 data_in =	-1068	;
#1000000 data_in =	-1093	;
#1000000 data_in =	-1110	;
#1000000 data_in =	-1135	;
#1000000 data_in =	-1152	;
#1000000 data_in =	-1178	;
#1000000 data_in =	-1194	;
#1000000 data_in =	-1220	;
#1000000 data_in =	-1253	;
#1000000 data_in =	-1279	;
#1000000 data_in =	-1321	;
#1000000 data_in =	-1354	;
#1000000 data_in =	-1396	;
#1000000 data_in =	-1439	;
#1000000 data_in =	-1489	;
#1000000 data_in =	-1531	;
#1000000 data_in =	-1573	;
#1000000 data_in =	-1615	;
#1000000 data_in =	-1649	;
#1000000 data_in =	-1683	;
#1000000 data_in =	-1708	;
#1000000 data_in =	-1716	;
#1000000 data_in =	-1725	;
#1000000 data_in =	-1725	;
#1000000 data_in =	-1708	;
#1000000 data_in =	-1683	;
#1000000 data_in =	-1641	;
#1000000 data_in =	-1590	;
#1000000 data_in =	-1531	;
#1000000 data_in =	-1464	;
#1000000 data_in =	-1388	;
#1000000 data_in =	-1312	;
#1000000 data_in =	-1220	;
#1000000 data_in =	-1127	;
#1000000 data_in =	-1043	;
#1000000 data_in =	-950	;
#1000000 data_in =	-866	;
#1000000 data_in =	-782	;
#1000000 data_in =	-706	;
#1000000 data_in =	-639	;
#1000000 data_in =	-580	;
#1000000 data_in =	-521	;
#1000000 data_in =	-470	;
#1000000 data_in =	-428	;
#1000000 data_in =	-386	;
#1000000 data_in =	-344	;
#1000000 data_in =	-310	;
#1000000 data_in =	-276	;
#1000000 data_in =	-243	;
#1000000 data_in =	-209	;
#1000000 data_in =	-175	;
#1000000 data_in =	-142	;
#1000000 data_in =	-108	;
#1000000 data_in =	-74	;
#1000000 data_in =	-49	;
#1000000 data_in =	-24	;
#1000000 data_in =	0	;
#1000000 data_in =	17	;
#1000000 data_in =	34	;
#1000000 data_in =	51	;
#1000000 data_in =	59	;
#1000000 data_in =	68	;
#1000000 data_in =	68	;
#1000000 data_in =	76	;
#1000000 data_in =	76	;
#1000000 data_in =	76	;
#1000000 data_in =	76	;
#1000000 data_in =	76	;
#1000000 data_in =	68	;
#1000000 data_in =	68	;
#1000000 data_in =	68	;
#1000000 data_in =	68	;
#1000000 data_in =	68	;
#1000000 data_in =	68	;
#1000000 data_in =	68	;
#1000000 data_in =	68	;
#1000000 data_in =	68	;
#1000000 data_in =	68	;
#1000000 data_in =	76	;
#1000000 data_in =	76	;
#1000000 data_in =	76	;
#1000000 data_in =	85	;
#1000000 data_in =	85	;
#1000000 data_in =	93	;
#1000000 data_in =	93	;
#1000000 data_in =	101	;
#1000000 data_in =	101	;
#1000000 data_in =	110	;
#1000000 data_in =	110	;
#1000000 data_in =	118	;
#1000000 data_in =	118	;
#1000000 data_in =	118	;
#1000000 data_in =	127	;
#1000000 data_in =	127	;
#1000000 data_in =	127	;
#1000000 data_in =	127	;
#1000000 data_in =	127	;
#1000000 data_in =	127	;
#1000000 data_in =	127	;
#1000000 data_in =	127	;
#1000000 data_in =	127	;
#1000000 data_in =	127	;
#1000000 data_in =	127	;
#1000000 data_in =	118	;
#1000000 data_in =	118	;
#1000000 data_in =	118	;
#1000000 data_in =	118	;
#1000000 data_in =	110	;
#1000000 data_in =	110	;
#1000000 data_in =	110	;
#1000000 data_in =	110	;
#1000000 data_in =	110	;
#1000000 data_in =	110	;
#1000000 data_in =	110	;
#1000000 data_in =	110	;
#1000000 data_in =	101	;
#1000000 data_in =	101	;
#1000000 data_in =	101	;
#1000000 data_in =	101	;
#1000000 data_in =	101	;
#1000000 data_in =	101	;
#1000000 data_in =	101	;
#1000000 data_in =	101	;
#1000000 data_in =	101	;
#1000000 data_in =	101	;
#1000000 data_in =	101	;
#1000000 data_in =	101	;
#1000000 data_in =	101	;
#1000000 data_in =	101	;
#1000000 data_in =	101	;
#1000000 data_in =	110	;
#1000000 data_in =	110	;
#1000000 data_in =	110	;
#1000000 data_in =	110	;
#1000000 data_in =	110	;
#1000000 data_in =	118	;
#1000000 data_in =	118	;
#1000000 data_in =	118	;
#1000000 data_in =	118	;
#1000000 data_in =	118	;
#1000000 data_in =	127	;
#1000000 data_in =	127	;
#1000000 data_in =	127	;
#1000000 data_in =	127	;
#1000000 data_in =	127	;
#1000000 data_in =	127	;
#1000000 data_in =	127	;
#1000000 data_in =	118	;
#1000000 data_in =	118	;
#1000000 data_in =	118	;
#1000000 data_in =	118	;
#1000000 data_in =	118	;
#1000000 data_in =	110	;
#1000000 data_in =	110	;
#1000000 data_in =	110	;
#1000000 data_in =	110	;
#1000000 data_in =	110	;
#1000000 data_in =	110	;
#1000000 data_in =	110	;
#1000000 data_in =	110	;
#1000000 data_in =	110	;
#1000000 data_in =	110	;
#1000000 data_in =	110	;
#1000000 data_in =	110	;
#1000000 data_in =	110	;
#1000000 data_in =	110	;
#1000000 data_in =	110	;
#1000000 data_in =	110	;
#1000000 data_in =	110	;
#1000000 data_in =	101	;
#1000000 data_in =	101	;
#1000000 data_in =	101	;
#1000000 data_in =	101	;
#1000000 data_in =	101	;
#1000000 data_in =	101	;
#1000000 data_in =	101	;
#1000000 data_in =	101	;
#1000000 data_in =	101	;
#1000000 data_in =	101	;
#1000000 data_in =	101	;
#1000000 data_in =	101	;
#1000000 data_in =	101	;
#1000000 data_in =	101	;
#1000000 data_in =	101	;
#1000000 data_in =	93	;
#1000000 data_in =	93	;
#1000000 data_in =	93	;
#1000000 data_in =	93	;
#1000000 data_in =	93	;
#1000000 data_in =	93	;
#1000000 data_in =	85	;
#1000000 data_in =	85	;
#1000000 data_in =	85	;
#1000000 data_in =	76	;
#1000000 data_in =	76	;
#1000000 data_in =	68	;
#1000000 data_in =	68	;
#1000000 data_in =	68	;
#1000000 data_in =	59	;
#1000000 data_in =	59	;
#1000000 data_in =	59	;
#1000000 data_in =	59	;
#1000000 data_in =	59	;
#1000000 data_in =	59	;
#1000000 data_in =	51	;
#1000000 data_in =	51	;
#1000000 data_in =	51	;
#1000000 data_in =	51	;
#1000000 data_in =	51	;
#1000000 data_in =	51	;
#1000000 data_in =	43	;
#1000000 data_in =	43	;
#1000000 data_in =	43	;
#1000000 data_in =	34	;
#1000000 data_in =	34	;
#1000000 data_in =	26	;
#1000000 data_in =	17	;
#1000000 data_in =	17	;
#1000000 data_in =	9	;
#1000000 data_in =	0	;
#1000000 data_in =	-7	;
#1000000 data_in =	-7	;
#1000000 data_in =	-15	;
#1000000 data_in =	-15	;
#1000000 data_in =	-24	;
#1000000 data_in =	-24	;
#1000000 data_in =	-32	;
#1000000 data_in =	-32	;
#1000000 data_in =	-41	;
#1000000 data_in =	-41	;
#1000000 data_in =	-41	;
#1000000 data_in =	-49	;
#1000000 data_in =	-49	;
#1000000 data_in =	-58	;
#1000000 data_in =	-58	;
#1000000 data_in =	-66	;
#1000000 data_in =	-74	;
#1000000 data_in =	-83	;
#1000000 data_in =	-83	;
#1000000 data_in =	-91	;
#1000000 data_in =	-100	;
#1000000 data_in =	-108	;
#1000000 data_in =	-116	;
#1000000 data_in =	-125	;
#1000000 data_in =	-133	;
#1000000 data_in =	-142	;
#1000000 data_in =	-150	;
#1000000 data_in =	-159	;
#1000000 data_in =	-167	;
#1000000 data_in =	-175	;
#1000000 data_in =	-184	;
#1000000 data_in =	-192	;
#1000000 data_in =	-201	;
#1000000 data_in =	-209	;
#1000000 data_in =	-218	;
#1000000 data_in =	-234	;
#1000000 data_in =	-243	;
#1000000 data_in =	-251	;
#1000000 data_in =	-260	;
#1000000 data_in =	-268	;
#1000000 data_in =	-285	;
#1000000 data_in =	-293	;
#1000000 data_in =	-302	;
#1000000 data_in =	-319	;
#1000000 data_in =	-327	;
#1000000 data_in =	-344	;
#1000000 data_in =	-361	;
#1000000 data_in =	-369	;
#1000000 data_in =	-386	;
#1000000 data_in =	-403	;
#1000000 data_in =	-420	;
#1000000 data_in =	-428	;
#1000000 data_in =	-445	;
#1000000 data_in =	-462	;
#1000000 data_in =	-470	;
#1000000 data_in =	-487	;
#1000000 data_in =	-504	;
#1000000 data_in =	-512	;
#1000000 data_in =	-529	;
#1000000 data_in =	-546	;
#1000000 data_in =	-563	;
#1000000 data_in =	-588	;
#1000000 data_in =	-605	;
#1000000 data_in =	-630	;
#1000000 data_in =	-647	;
#1000000 data_in =	-672	;
#1000000 data_in =	-698	;
#1000000 data_in =	-714	;
#1000000 data_in =	-740	;
#1000000 data_in =	-765	;
#1000000 data_in =	-790	;
#1000000 data_in =	-807	;
#1000000 data_in =	-832	;
#1000000 data_in =	-858	;
#1000000 data_in =	-874	;
#1000000 data_in =	-891	;
#1000000 data_in =	-908	;
#1000000 data_in =	-933	;
#1000000 data_in =	-950	;
#1000000 data_in =	-967	;
#1000000 data_in =	-984	;
#1000000 data_in =	-1001	;
#1000000 data_in =	-1018	;
#1000000 data_in =	-1034	;
#1000000 data_in =	-1060	;
#1000000 data_in =	-1076	;
#1000000 data_in =	-1093	;
#1000000 data_in =	-1119	;
#1000000 data_in =	-1135	;
#1000000 data_in =	-1161	;
#1000000 data_in =	-1186	;
#1000000 data_in =	-1203	;
#1000000 data_in =	-1228	;
#1000000 data_in =	-1245	;
#1000000 data_in =	-1270	;
#1000000 data_in =	-1287	;
#1000000 data_in =	-1304	;
#1000000 data_in =	-1329	;
#1000000 data_in =	-1346	;
#1000000 data_in =	-1363	;
#1000000 data_in =	-1371	;
#1000000 data_in =	-1388	;
#1000000 data_in =	-1405	;
#1000000 data_in =	-1413	;
#1000000 data_in =	-1430	;
#1000000 data_in =	-1439	;
#1000000 data_in =	-1447	;
#1000000 data_in =	-1455	;
#1000000 data_in =	-1472	;
#1000000 data_in =	-1481	;
#1000000 data_in =	-1489	;
#1000000 data_in =	-1498	;
#1000000 data_in =	-1506	;
#1000000 data_in =	-1514	;
#1000000 data_in =	-1523	;
#1000000 data_in =	-1531	;
#1000000 data_in =	-1540	;
#1000000 data_in =	-1548	;
#1000000 data_in =	-1556	;
#1000000 data_in =	-1556	;
#1000000 data_in =	-1565	;
#1000000 data_in =	-1565	;
#1000000 data_in =	-1565	;
#1000000 data_in =	-1565	;
#1000000 data_in =	-1565	;
#1000000 data_in =	-1565	;
#1000000 data_in =	-1565	;
#1000000 data_in =	-1565	;
#1000000 data_in =	-1565	;
#1000000 data_in =	-1556	;
#1000000 data_in =	-1556	;
#1000000 data_in =	-1556	;
#1000000 data_in =	-1548	;
#1000000 data_in =	-1540	;
#1000000 data_in =	-1540	;
#1000000 data_in =	-1531	;
#1000000 data_in =	-1523	;
#1000000 data_in =	-1506	;
#1000000 data_in =	-1498	;
#1000000 data_in =	-1489	;
#1000000 data_in =	-1472	;
#1000000 data_in =	-1455	;
#1000000 data_in =	-1439	;
#1000000 data_in =	-1413	;
#1000000 data_in =	-1396	;
#1000000 data_in =	-1371	;
#1000000 data_in =	-1354	;
#1000000 data_in =	-1329	;
#1000000 data_in =	-1304	;
#1000000 data_in =	-1279	;
#1000000 data_in =	-1253	;
#1000000 data_in =	-1220	;
#1000000 data_in =	-1194	;
#1000000 data_in =	-1169	;
#1000000 data_in =	-1144	;
#1000000 data_in =	-1110	;
#1000000 data_in =	-1085	;
#1000000 data_in =	-1060	;
#1000000 data_in =	-1026	;
#1000000 data_in =	-1001	;
#1000000 data_in =	-975	;
#1000000 data_in =	-942	;
#1000000 data_in =	-916	;
#1000000 data_in =	-891	;
#1000000 data_in =	-866	;
#1000000 data_in =	-841	;
#1000000 data_in =	-815	;
#1000000 data_in =	-799	;
#1000000 data_in =	-773	;
#1000000 data_in =	-748	;
#1000000 data_in =	-723	;
#1000000 data_in =	-698	;
#1000000 data_in =	-664	;
#1000000 data_in =	-639	;
#1000000 data_in =	-613	;
#1000000 data_in =	-580	;
#1000000 data_in =	-554	;
#1000000 data_in =	-521	;
#1000000 data_in =	-495	;
#1000000 data_in =	-470	;
#1000000 data_in =	-445	;
#1000000 data_in =	-420	;
#1000000 data_in =	-394	;
#1000000 data_in =	-378	;
#1000000 data_in =	-352	;
#1000000 data_in =	-335	;
#1000000 data_in =	-319	;
#1000000 data_in =	-302	;
#1000000 data_in =	-285	;
#1000000 data_in =	-276	;
#1000000 data_in =	-260	;
#1000000 data_in =	-243	;
#1000000 data_in =	-226	;
#1000000 data_in =	-218	;
#1000000 data_in =	-201	;
#1000000 data_in =	-184	;
#1000000 data_in =	-175	;
#1000000 data_in =	-159	;
#1000000 data_in =	-142	;
#1000000 data_in =	-133	;
#1000000 data_in =	-125	;
#1000000 data_in =	-108	;
#1000000 data_in =	-100	;
#1000000 data_in =	-91	;
#1000000 data_in =	-83	;
#1000000 data_in =	-74	;
#1000000 data_in =	-74	;
#1000000 data_in =	-66	;
#1000000 data_in =	-58	;
#1000000 data_in =	-49	;
#1000000 data_in =	-49	;
#1000000 data_in =	-41	;
#1000000 data_in =	-32	;
#1000000 data_in =	-24	;
#1000000 data_in =	-24	;
#1000000 data_in =	-15	;
#1000000 data_in =	-7	;
#1000000 data_in =	-7	;
#1000000 data_in =	0	;
#1000000 data_in =	0	;
#1000000 data_in =	9	;
#1000000 data_in =	9	;
#1000000 data_in =	17	;
#1000000 data_in =	17	;
#1000000 data_in =	26	;
#1000000 data_in =	26	;
#1000000 data_in =	34	;
#1000000 data_in =	34	;
#1000000 data_in =	34	;
#1000000 data_in =	43	;
#1000000 data_in =	43	;
#1000000 data_in =	51	;
#1000000 data_in =	51	;
#1000000 data_in =	59	;
#1000000 data_in =	59	;
#1000000 data_in =	68	;
#1000000 data_in =	68	;
#1000000 data_in =	76	;
#1000000 data_in =	76	;
#1000000 data_in =	76	;
#1000000 data_in =	85	;
#1000000 data_in =	85	;
#1000000 data_in =	93	;
#1000000 data_in =	93	;
#1000000 data_in =	93	;
#1000000 data_in =	101	;
#1000000 data_in =	101	;
#1000000 data_in =	101	;
#1000000 data_in =	101	;
#1000000 data_in =	101	;
#1000000 data_in =	110	;
#1000000 data_in =	110	;
#1000000 data_in =	110	;
#1000000 data_in =	110	;
#1000000 data_in =	110	;
#1000000 data_in =	118	;
#1000000 data_in =	118	;
#1000000 data_in =	118	;
#1000000 data_in =	118	;
#1000000 data_in =	118	;
#1000000 data_in =	127	;
#1000000 data_in =	127	;
#1000000 data_in =	127	;
#1000000 data_in =	127	;
#1000000 data_in =	127	;
#1000000 data_in =	135	;
#1000000 data_in =	135	;
#1050000 data_in =	1	;
#1000000 data_in = 	30	;



end

endmodule


