`timescale 1ns / 100ps
`include "parameter.v"

module waveletl5 (q_peak_ref,q_peak_pos_ref,s_peak_ref,s_peak_pos_ref,p_begin,
p_end,p_peak,p_peak_pos,t_begin,t_end,t_peak,t_peak_pos,
start_qrs_fin_2,end_qrs_fin_2,r_peak_pos_ref,
ecg0,ecg1,ecg2,ecg3,ecg4,ecg5,ecg6,ecg7,ecg8,ecg9,ecg10,ecg11,ecg12,ecg13,ecg14,ecg15,ecg16,ecg17,ecg18,ecg19,ecg20,ecg21,ecg22,ecg23,ecg24,ecg25,ecg26,ecg27,ecg28,ecg29,ecg30,ecg31,ecg32,ecg33,ecg34,ecg35,ecg36,ecg37,ecg38,ecg39,ecg40,ecg41,ecg42,ecg43,ecg44,ecg45,ecg46,ecg47,ecg48,ecg49,ecg50,ecg51,ecg52,ecg53,ecg54,ecg55,ecg56,ecg57,ecg58,ecg59,ecg60,ecg61,ecg62,ecg63,ecg64,ecg65,ecg66,ecg67,ecg68,ecg69,ecg70,ecg71,ecg72,ecg73,ecg74,ecg75,ecg76,ecg77,ecg78,ecg79,ecg80,ecg81,ecg82,ecg83,ecg84,ecg85,ecg86,ecg87,ecg88,ecg89,ecg90,ecg91,ecg92,ecg93,ecg94,ecg95,ecg96,ecg97,ecg98,ecg99,ecg100,ecg101,ecg102,ecg103,ecg104,ecg105,ecg106,ecg107,ecg108,ecg109,ecg110,ecg111,ecg112,ecg113,ecg114,ecg115,ecg116,ecg117,ecg118,ecg119,ecg120,ecg121,ecg122,ecg123,ecg124,ecg125,ecg126,ecg127,ecg128,ecg129,ecg130,ecg131,ecg132,ecg133,ecg134,ecg135,ecg136,ecg137,ecg138,ecg139,ecg140,ecg141,ecg142,ecg143,ecg144,ecg145,ecg146,ecg147,ecg148,ecg149,ecg150,ecg151,ecg152,ecg153,ecg154,ecg155,ecg156,ecg157,ecg158,ecg159,ecg160,ecg161,ecg162,ecg163,ecg164,ecg165,ecg166,ecg167,ecg168,ecg169,ecg170,ecg171,ecg172,ecg173,ecg174,ecg175,ecg176,ecg177,ecg178,ecg179,ecg180,ecg181,ecg182,ecg183,ecg184,ecg185,ecg186,ecg187,ecg188,ecg189,ecg190,ecg191,ecg192,ecg193,ecg194,ecg195,ecg196,ecg197,ecg198,ecg199,ecg200,ecg201,ecg202,ecg203,ecg204,ecg205,ecg206,ecg207,ecg208,ecg209,ecg210,ecg211,ecg212,ecg213,ecg214,ecg215,ecg216,ecg217,ecg218,ecg219,ecg220,ecg221,ecg222,ecg223,ecg224,ecg225,ecg226,ecg227,ecg228,ecg229,ecg230,ecg231,ecg232,ecg233,ecg234,ecg235,ecg236,ecg237,ecg238,ecg239,ecg240,ecg241,ecg242,ecg243,ecg244,ecg245,ecg246,ecg247,ecg248,ecg249,ecg250,ecg251,ecg252,ecg253,ecg254,ecg255,ecg256,ecg257,ecg258,ecg259,ecg260,ecg261,ecg262,ecg263,ecg264,ecg265,ecg266,ecg267,ecg268,ecg269,ecg270,ecg271,ecg272,ecg273,ecg274,ecg275,ecg276,ecg277,ecg278,ecg279,ecg280,ecg281,ecg282,ecg283,ecg284,ecg285,ecg286,ecg287,ecg288,ecg289,ecg290,ecg291,ecg292,ecg293,ecg294,ecg295,ecg296,ecg297,ecg298,ecg299,ecg300,ecg301,ecg302,ecg303,ecg304,ecg305,ecg306,ecg307,ecg308,ecg309,ecg310,ecg311,ecg312,ecg313,ecg314,ecg315,ecg316,ecg317,ecg318,ecg319,ecg320,ecg321,ecg322,ecg323,ecg324,ecg325,ecg326,ecg327,ecg328,ecg329,ecg330,ecg331,ecg332,ecg333,ecg334,ecg335,ecg336,ecg337,ecg338,ecg339,ecg340,ecg341,ecg342,ecg343,ecg344,ecg345,ecg346,ecg347,ecg348,ecg349,ecg350,ecg351,ecg352,ecg353,ecg354,ecg355,ecg356,ecg357,ecg358,ecg359,ecg360,ecg361,ecg362,ecg363,ecg364,ecg365,ecg366,ecg367,ecg368,ecg369,ecg370,ecg371,ecg372,ecg373,ecg374,ecg375,ecg376,ecg377,ecg378,ecg379,ecg380,ecg381,ecg382,ecg383,ecg384,ecg385,ecg386,ecg387,ecg388,ecg389,ecg390,ecg391,ecg392,ecg393,ecg394,ecg395,ecg396,ecg397,ecg398,ecg399,ecg400,ecg401,ecg402,ecg403,ecg404,ecg405,ecg406,ecg407,ecg408,ecg409,ecg410,ecg411,ecg412,ecg413,ecg414,ecg415,ecg416,ecg417,ecg418,ecg419,ecg420,ecg421,ecg422,ecg423,ecg424,ecg425,ecg426,ecg427,ecg428,ecg429,ecg430,ecg431,ecg432,ecg433,ecg434,ecg435,ecg436,ecg437,ecg438,ecg439,ecg440,ecg441,ecg442,ecg443,ecg444,ecg445,ecg446,ecg447,ecg448,ecg449,ecg450,ecg451,ecg452,ecg453,ecg454,ecg455,ecg456,ecg457,ecg458,ecg459,ecg460,ecg461,ecg462,ecg463,ecg464,ecg465,ecg466,ecg467,ecg468,ecg469,ecg470,ecg471,ecg472,ecg473,ecg474,ecg475,ecg476,ecg477,ecg478,ecg479,ecg480,ecg481,ecg482,ecg483,ecg484,ecg485,ecg486,ecg487,ecg488,ecg489,ecg490,ecg491,ecg492,ecg493,ecg494,ecg495,ecg496,ecg497,ecg498,ecg499,ecg500,ecg501,ecg502,ecg503,ecg504,ecg505,ecg506,ecg507,ecg508,ecg509,ecg510,ecg511,ecg512,ecg513,ecg514,ecg515,ecg516,ecg517,ecg518,ecg519,ecg520,ecg521,ecg522,ecg523,ecg524,ecg525,ecg526,ecg527,ecg528,ecg529,ecg530,ecg531,ecg532,ecg533,ecg534,ecg535,ecg536,ecg537,ecg538,ecg539,ecg540,ecg541,ecg542,ecg543,ecg544,ecg545,ecg546,ecg547,ecg548,ecg549,ecg550,ecg551,ecg552,ecg553,ecg554,ecg555,ecg556,ecg557,ecg558,ecg559,ecg560,ecg561,ecg562,ecg563,ecg564,ecg565,ecg566,ecg567,ecg568,ecg569,ecg570,ecg571,ecg572,ecg573,ecg574,ecg575,ecg576,ecg577,ecg578,ecg579,ecg580,ecg581,ecg582,ecg583,ecg584,ecg585,ecg586,ecg587,ecg588,ecg589,ecg590,ecg591,ecg592,ecg593,ecg594,ecg595,ecg596,ecg597,ecg598,ecg599,
ecg600,ecg601,ecg602,ecg603,ecg604,ecg605,ecg606,ecg607,ecg608,ecg609,ecg610,ecg611,ecg612,ecg613,ecg614,ecg615,ecg616,ecg617,ecg618,ecg619,ecg620,ecg621,ecg622,ecg623,ecg624,ecg625,ecg626,ecg627,ecg628,ecg629,ecg630,ecg631,ecg632,ecg633,ecg634,ecg635,ecg636,ecg637,ecg638,ecg639,ecg640,ecg641,ecg642,ecg643,ecg644,ecg645,ecg646,ecg647,ecg648,ecg649,ecg650,ecg651,ecg652,ecg653,ecg654,ecg655,ecg656,ecg657,ecg658,ecg659,ecg660,ecg661,ecg662,ecg663,ecg664,ecg665,ecg666,ecg667,ecg668,ecg669,ecg670,ecg671,ecg672,ecg673,ecg674,ecg675,ecg676,ecg677,ecg678,ecg679,ecg680,ecg681,ecg682,ecg683,ecg684,ecg685,ecg686,ecg687,ecg688,ecg689,ecg690,ecg691,ecg692,ecg693,ecg694,ecg695,ecg696,ecg697,ecg698,ecg699,ecg700,ecg701,ecg702,ecg703,ecg704,ecg705,ecg706,ecg707,ecg708,ecg709,ecg710,ecg711,ecg712,ecg713,ecg714,ecg715,ecg716,ecg717,ecg718,ecg719,ecg720,ecg721,ecg722,ecg723,ecg724,ecg725,ecg726,ecg727,ecg728,ecg729,ecg730,ecg731,ecg732,ecg733,ecg734,ecg735,ecg736,ecg737,ecg738,ecg739,ecg740,ecg741,ecg742,ecg743,ecg744,ecg745,ecg746,ecg747,ecg748,ecg749,ecg750,ecg751,ecg752,ecg753,ecg754,ecg755,ecg756,ecg757,ecg758,ecg759,ecg760,ecg761,ecg762,ecg763,ecg764,ecg765,ecg766,ecg767,ecg768,ecg769,ecg770,ecg771,ecg772,ecg773,ecg774,ecg775,ecg776,ecg777,ecg778,ecg779,ecg780,ecg781,ecg782,ecg783,ecg784,ecg785,ecg786,ecg787,ecg788,ecg789,ecg790,ecg791,ecg792,ecg793,ecg794,ecg795,ecg796,ecg797,ecg798,ecg799,data_in,clk,nReset);

output signed [15:0] q_peak_ref,q_peak_pos_ref,s_peak_ref,s_peak_pos_ref,p_begin,p_end,p_peak,p_peak_pos,t_begin,t_end,t_peak,t_peak_pos; 

input signed [15:0] start_qrs_fin_2,end_qrs_fin_2,r_peak_pos_ref,
ecg0,ecg1,ecg2,ecg3,ecg4,ecg5,ecg6,ecg7,ecg8,ecg9,ecg10,ecg11,ecg12,ecg13,ecg14,ecg15,ecg16,ecg17,ecg18,ecg19,ecg20,ecg21,ecg22,ecg23,ecg24,ecg25,ecg26,ecg27,ecg28,ecg29,ecg30,ecg31,ecg32,ecg33,ecg34,ecg35,ecg36,ecg37,ecg38,ecg39,ecg40,ecg41,ecg42,ecg43,ecg44,ecg45,ecg46,ecg47,ecg48,ecg49,ecg50,ecg51,ecg52,ecg53,ecg54,ecg55,ecg56,ecg57,ecg58,ecg59,ecg60,ecg61,ecg62,ecg63,ecg64,ecg65,ecg66,ecg67,ecg68,ecg69,ecg70,ecg71,ecg72,ecg73,ecg74,ecg75,ecg76,ecg77,ecg78,ecg79,ecg80,ecg81,ecg82,ecg83,ecg84,ecg85,ecg86,ecg87,ecg88,ecg89,ecg90,ecg91,ecg92,ecg93,ecg94,ecg95,ecg96,ecg97,ecg98,ecg99,ecg100,ecg101,ecg102,ecg103,ecg104,ecg105,ecg106,ecg107,ecg108,ecg109,ecg110,ecg111,ecg112,ecg113,ecg114,ecg115,ecg116,ecg117,ecg118,ecg119,ecg120,ecg121,ecg122,ecg123,ecg124,ecg125,ecg126,ecg127,ecg128,ecg129,ecg130,ecg131,ecg132,ecg133,ecg134,ecg135,ecg136,ecg137,ecg138,ecg139,ecg140,ecg141,ecg142,ecg143,ecg144,ecg145,ecg146,ecg147,ecg148,ecg149,ecg150,ecg151,ecg152,ecg153,ecg154,ecg155,ecg156,ecg157,ecg158,ecg159,ecg160,ecg161,ecg162,ecg163,ecg164,ecg165,ecg166,ecg167,ecg168,ecg169,ecg170,ecg171,ecg172,ecg173,ecg174,ecg175,ecg176,ecg177,ecg178,ecg179,ecg180,ecg181,ecg182,ecg183,ecg184,ecg185,ecg186,ecg187,ecg188,ecg189,ecg190,ecg191,ecg192,ecg193,ecg194,ecg195,ecg196,ecg197,ecg198,ecg199,ecg200,ecg201,ecg202,ecg203,ecg204,ecg205,ecg206,ecg207,ecg208,ecg209,ecg210,ecg211,ecg212,ecg213,ecg214,ecg215,ecg216,ecg217,ecg218,ecg219,ecg220,ecg221,ecg222,ecg223,ecg224,ecg225,ecg226,ecg227,ecg228,ecg229,ecg230,ecg231,ecg232,ecg233,ecg234,ecg235,ecg236,ecg237,ecg238,ecg239,ecg240,ecg241,ecg242,ecg243,ecg244,ecg245,ecg246,ecg247,ecg248,ecg249,ecg250,ecg251,ecg252,ecg253,ecg254,ecg255,ecg256,ecg257,ecg258,ecg259,ecg260,ecg261,ecg262,ecg263,ecg264,ecg265,ecg266,ecg267,ecg268,ecg269,ecg270,ecg271,ecg272,ecg273,ecg274,ecg275,ecg276,ecg277,ecg278,ecg279,ecg280,ecg281,ecg282,ecg283,ecg284,ecg285,ecg286,ecg287,ecg288,ecg289,ecg290,ecg291,ecg292,ecg293,ecg294,ecg295,ecg296,ecg297,ecg298,ecg299,ecg300,ecg301,ecg302,ecg303,ecg304,ecg305,ecg306,ecg307,ecg308,ecg309,ecg310,ecg311,ecg312,ecg313,ecg314,ecg315,ecg316,ecg317,ecg318,ecg319,ecg320,ecg321,ecg322,ecg323,ecg324,ecg325,ecg326,ecg327,ecg328,ecg329,ecg330,ecg331,ecg332,ecg333,ecg334,ecg335,ecg336,ecg337,ecg338,ecg339,ecg340,ecg341,ecg342,ecg343,ecg344,ecg345,ecg346,ecg347,ecg348,ecg349,ecg350,ecg351,ecg352,ecg353,ecg354,ecg355,ecg356,ecg357,ecg358,ecg359,ecg360,ecg361,ecg362,ecg363,ecg364,ecg365,ecg366,ecg367,ecg368,ecg369,ecg370,ecg371,ecg372,ecg373,ecg374,ecg375,ecg376,ecg377,ecg378,ecg379,ecg380,ecg381,ecg382,ecg383,ecg384,ecg385,ecg386,ecg387,ecg388,ecg389,ecg390,ecg391,ecg392,ecg393,ecg394,ecg395,ecg396,ecg397,ecg398,ecg399,ecg400,ecg401,ecg402,ecg403,ecg404,ecg405,ecg406,ecg407,ecg408,ecg409,ecg410,ecg411,ecg412,ecg413,ecg414,ecg415,ecg416,ecg417,ecg418,ecg419,ecg420,ecg421,ecg422,ecg423,ecg424,ecg425,ecg426,ecg427,ecg428,ecg429,ecg430,ecg431,ecg432,ecg433,ecg434,ecg435,ecg436,ecg437,ecg438,ecg439,ecg440,ecg441,ecg442,ecg443,ecg444,ecg445,ecg446,ecg447,ecg448,ecg449,ecg450,ecg451,ecg452,ecg453,ecg454,ecg455,ecg456,ecg457,ecg458,ecg459,ecg460,ecg461,ecg462,ecg463,ecg464,ecg465,ecg466,ecg467,ecg468,ecg469,ecg470,ecg471,ecg472,ecg473,ecg474,ecg475,ecg476,ecg477,ecg478,ecg479,ecg480,ecg481,ecg482,ecg483,ecg484,ecg485,ecg486,ecg487,ecg488,ecg489,ecg490,ecg491,ecg492,ecg493,ecg494,ecg495,ecg496,ecg497,ecg498,ecg499,ecg500,ecg501,ecg502,ecg503,ecg504,ecg505,ecg506,ecg507,ecg508,ecg509,ecg510,ecg511,ecg512,ecg513,ecg514,ecg515,ecg516,ecg517,ecg518,ecg519,ecg520,ecg521,ecg522,ecg523,ecg524,ecg525,ecg526,ecg527,ecg528,ecg529,ecg530,ecg531,ecg532,ecg533,ecg534,ecg535,ecg536,ecg537,ecg538,ecg539,ecg540,ecg541,ecg542,ecg543,ecg544,ecg545,ecg546,ecg547,ecg548,ecg549,ecg550,ecg551,ecg552,ecg553,ecg554,ecg555,ecg556,ecg557,ecg558,ecg559,ecg560,ecg561,ecg562,ecg563,ecg564,ecg565,ecg566,ecg567,ecg568,ecg569,ecg570,ecg571,ecg572,ecg573,ecg574,ecg575,ecg576,ecg577,ecg578,ecg579,ecg580,ecg581,ecg582,ecg583,ecg584,ecg585,ecg586,ecg587,ecg588,ecg589,ecg590,ecg591,ecg592,ecg593,ecg594,ecg595,ecg596,ecg597,ecg598,ecg599,
ecg600,ecg601,ecg602,ecg603,ecg604,ecg605,ecg606,ecg607,ecg608,ecg609,ecg610,ecg611,ecg612,ecg613,ecg614,ecg615,ecg616,ecg617,ecg618,ecg619,ecg620,ecg621,ecg622,ecg623,ecg624,ecg625,ecg626,ecg627,ecg628,ecg629,ecg630,ecg631,ecg632,ecg633,ecg634,ecg635,ecg636,ecg637,ecg638,ecg639,ecg640,ecg641,ecg642,ecg643,ecg644,ecg645,ecg646,ecg647,ecg648,ecg649,ecg650,ecg651,ecg652,ecg653,ecg654,ecg655,ecg656,ecg657,ecg658,ecg659,ecg660,ecg661,ecg662,ecg663,ecg664,ecg665,ecg666,ecg667,ecg668,ecg669,ecg670,ecg671,ecg672,ecg673,ecg674,ecg675,ecg676,ecg677,ecg678,ecg679,ecg680,ecg681,ecg682,ecg683,ecg684,ecg685,ecg686,ecg687,ecg688,ecg689,ecg690,ecg691,ecg692,ecg693,ecg694,ecg695,ecg696,ecg697,ecg698,ecg699,ecg700,ecg701,ecg702,ecg703,ecg704,ecg705,ecg706,ecg707,ecg708,ecg709,ecg710,ecg711,ecg712,ecg713,ecg714,ecg715,ecg716,ecg717,ecg718,ecg719,ecg720,ecg721,ecg722,ecg723,ecg724,ecg725,ecg726,ecg727,ecg728,ecg729,ecg730,ecg731,ecg732,ecg733,ecg734,ecg735,ecg736,ecg737,ecg738,ecg739,ecg740,ecg741,ecg742,ecg743,ecg744,ecg745,ecg746,ecg747,ecg748,ecg749,ecg750,ecg751,ecg752,ecg753,ecg754,ecg755,ecg756,ecg757,ecg758,ecg759,ecg760,ecg761,ecg762,ecg763,ecg764,ecg765,ecg766,ecg767,ecg768,ecg769,ecg770,ecg771,ecg772,ecg773,ecg774,ecg775,ecg776,ecg777,ecg778,ecg779,ecg780,ecg781,ecg782,ecg783,ecg784,ecg785,ecg786,ecg787,ecg788,ecg789,ecg790,ecg791,ecg792,ecg793,ecg794,ecg795,ecg796,ecg797,ecg798,ecg799;

input [15:0] data_in;

input clk, nReset;
wire clk, nReset;

wire [5:0] count1_l5,count2_l5;

wire signed [15:0] p1maxp,p1minp,p2maxp,p2minp,t1maxp,t1minp;

wire array_2,p1_cD_full,p2_cD_full,t_cD_full,p_zero;

level5arch l5arch(p_begin,p_end,p1maxp,p1minp,p2maxp,p2minp,t_begin,t_end,t1maxp,
t1minp,array_2,p1_cD_full,p2_cD_full,t_cD_full,p_zero,count1_l5,
count2_l5,start_qrs_fin_2,end_qrs_fin_2,data_in,clk,nReset);

ecg_signal_maxmin ecg_mxmn(q_peak_ref,q_peak_pos_ref,s_peak_ref,s_peak_pos_ref,p_peak,p_peak_pos,p_begin,p_end,t_peak,t_peak_pos,t_begin,t_end,array_2,
p1_cD_full,p2_cD_full,t_cD_full,p_zero,p1maxp,p1minp,
p2maxp,p2minp,t1maxp,t1minp,start_qrs_fin_2,end_qrs_fin_2,
r_peak_pos_ref,count1_l5,count2_l5,
ecg0,ecg1,ecg2,ecg3,ecg4,ecg5,ecg6,ecg7,ecg8,ecg9,
ecg10,ecg11,ecg12,ecg13,ecg14,ecg15,ecg16,ecg17,ecg18,ecg19,
ecg20,ecg21,ecg22,ecg23,ecg24,ecg25,ecg26,ecg27,ecg28,ecg29,ecg30,ecg31,ecg32,ecg33,ecg34,ecg35,ecg36,ecg37,ecg38,ecg39,ecg40,ecg41,ecg42,ecg43,ecg44,ecg45,ecg46,ecg47,ecg48,ecg49,ecg50,ecg51,ecg52,ecg53,ecg54,ecg55,ecg56,ecg57,ecg58,ecg59,ecg60,ecg61,ecg62,ecg63,ecg64,ecg65,ecg66,ecg67,ecg68,ecg69,ecg70,ecg71,ecg72,ecg73,ecg74,ecg75,ecg76,ecg77,ecg78,ecg79,ecg80,ecg81,ecg82,ecg83,ecg84,ecg85,ecg86,ecg87,ecg88,ecg89,ecg90,ecg91,ecg92,ecg93,ecg94,ecg95,ecg96,ecg97,ecg98,ecg99,ecg100,ecg101,ecg102,ecg103,ecg104,ecg105,ecg106,ecg107,ecg108,ecg109,ecg110,ecg111,ecg112,ecg113,ecg114,ecg115,ecg116,ecg117,ecg118,ecg119,ecg120,ecg121,ecg122,ecg123,ecg124,ecg125,ecg126,ecg127,ecg128,ecg129,ecg130,ecg131,ecg132,ecg133,ecg134,ecg135,ecg136,ecg137,ecg138,ecg139,ecg140,ecg141,ecg142,ecg143,ecg144,ecg145,ecg146,ecg147,ecg148,ecg149,ecg150,ecg151,ecg152,ecg153,ecg154,ecg155,ecg156,ecg157,ecg158,ecg159,ecg160,ecg161,ecg162,ecg163,ecg164,ecg165,ecg166,ecg167,ecg168,ecg169,ecg170,ecg171,ecg172,ecg173,ecg174,ecg175,ecg176,ecg177,ecg178,ecg179,ecg180,ecg181,ecg182,ecg183,ecg184,ecg185,ecg186,ecg187,ecg188,ecg189,ecg190,ecg191,ecg192,ecg193,ecg194,ecg195,ecg196,ecg197,ecg198,ecg199,ecg200,ecg201,ecg202,ecg203,ecg204,ecg205,ecg206,ecg207,ecg208,ecg209,ecg210,ecg211,ecg212,ecg213,ecg214,ecg215,ecg216,ecg217,ecg218,ecg219,ecg220,ecg221,ecg222,ecg223,ecg224,ecg225,ecg226,ecg227,ecg228,ecg229,ecg230,ecg231,ecg232,ecg233,ecg234,ecg235,ecg236,ecg237,ecg238,ecg239,ecg240,ecg241,ecg242,ecg243,ecg244,ecg245,ecg246,ecg247,ecg248,ecg249,ecg250,ecg251,ecg252,ecg253,ecg254,ecg255,ecg256,ecg257,ecg258,ecg259,ecg260,ecg261,ecg262,ecg263,ecg264,ecg265,ecg266,ecg267,ecg268,ecg269,ecg270,ecg271,ecg272,ecg273,ecg274,ecg275,ecg276,ecg277,ecg278,ecg279,ecg280,ecg281,ecg282,ecg283,ecg284,ecg285,ecg286,ecg287,ecg288,ecg289,ecg290,ecg291,ecg292,ecg293,ecg294,ecg295,ecg296,ecg297,ecg298,ecg299,ecg300,ecg301,ecg302,ecg303,ecg304,ecg305,ecg306,ecg307,ecg308,ecg309,ecg310,ecg311,ecg312,ecg313,ecg314,ecg315,ecg316,ecg317,ecg318,ecg319,ecg320,ecg321,ecg322,ecg323,ecg324,ecg325,ecg326,ecg327,ecg328,ecg329,ecg330,ecg331,ecg332,ecg333,ecg334,ecg335,ecg336,ecg337,ecg338,ecg339,ecg340,ecg341,ecg342,ecg343,ecg344,ecg345,ecg346,ecg347,ecg348,ecg349,ecg350,ecg351,ecg352,ecg353,ecg354,ecg355,ecg356,ecg357,ecg358,ecg359,ecg360,ecg361,ecg362,ecg363,ecg364,ecg365,ecg366,ecg367,ecg368,ecg369,ecg370,ecg371,ecg372,ecg373,ecg374,ecg375,ecg376,ecg377,ecg378,ecg379,ecg380,ecg381,ecg382,ecg383,ecg384,ecg385,ecg386,ecg387,ecg388,ecg389,ecg390,ecg391,ecg392,ecg393,ecg394,ecg395,ecg396,ecg397,ecg398,ecg399,ecg400,ecg401,ecg402,ecg403,ecg404,ecg405,ecg406,ecg407,ecg408,ecg409,ecg410,ecg411,ecg412,ecg413,ecg414,ecg415,ecg416,ecg417,ecg418,ecg419,ecg420,ecg421,ecg422,ecg423,ecg424,ecg425,ecg426,ecg427,ecg428,ecg429,ecg430,ecg431,ecg432,ecg433,ecg434,ecg435,ecg436,ecg437,ecg438,ecg439,ecg440,ecg441,ecg442,ecg443,ecg444,ecg445,ecg446,ecg447,ecg448,ecg449,ecg450,ecg451,ecg452,ecg453,ecg454,ecg455,ecg456,ecg457,ecg458,ecg459,ecg460,ecg461,ecg462,ecg463,ecg464,ecg465,ecg466,ecg467,ecg468,ecg469,ecg470,ecg471,ecg472,ecg473,ecg474,ecg475,ecg476,ecg477,ecg478,ecg479,ecg480,ecg481,ecg482,ecg483,ecg484,ecg485,ecg486,ecg487,ecg488,ecg489,ecg490,ecg491,ecg492,ecg493,ecg494,ecg495,ecg496,ecg497,ecg498,ecg499,ecg500,ecg501,ecg502,ecg503,ecg504,ecg505,ecg506,ecg507,ecg508,ecg509,ecg510,ecg511,ecg512,ecg513,ecg514,ecg515,ecg516,ecg517,ecg518,ecg519,ecg520,ecg521,ecg522,ecg523,ecg524,ecg525,ecg526,ecg527,ecg528,ecg529,ecg530,ecg531,ecg532,ecg533,ecg534,ecg535,ecg536,ecg537,ecg538,ecg539,ecg540,ecg541,ecg542,ecg543,ecg544,ecg545,ecg546,ecg547,ecg548,ecg549,ecg550,ecg551,ecg552,ecg553,ecg554,ecg555,ecg556,ecg557,ecg558,ecg559,ecg560,ecg561,ecg562,ecg563,ecg564,ecg565,ecg566,ecg567,ecg568,ecg569,ecg570,ecg571,ecg572,ecg573,ecg574,ecg575,ecg576,ecg577,ecg578,ecg579,ecg580,ecg581,ecg582,ecg583,ecg584,ecg585,ecg586,ecg587,ecg588,ecg589,ecg590,ecg591,ecg592,ecg593,ecg594,ecg595,ecg596,ecg597,ecg598,ecg599,
ecg600,ecg601,ecg602,ecg603,ecg604,ecg605,ecg606,ecg607,ecg608,ecg609,ecg610,ecg611,ecg612,ecg613,ecg614,ecg615,ecg616,ecg617,ecg618,ecg619,ecg620,ecg621,ecg622,ecg623,ecg624,ecg625,ecg626,ecg627,ecg628,ecg629,ecg630,ecg631,ecg632,ecg633,ecg634,ecg635,ecg636,ecg637,ecg638,ecg639,ecg640,ecg641,ecg642,ecg643,ecg644,ecg645,ecg646,ecg647,ecg648,ecg649,ecg650,ecg651,ecg652,ecg653,ecg654,ecg655,ecg656,ecg657,ecg658,ecg659,ecg660,ecg661,ecg662,ecg663,ecg664,ecg665,ecg666,ecg667,ecg668,ecg669,ecg670,ecg671,ecg672,ecg673,ecg674,ecg675,ecg676,ecg677,ecg678,ecg679,ecg680,ecg681,ecg682,ecg683,ecg684,ecg685,ecg686,ecg687,ecg688,ecg689,ecg690,ecg691,ecg692,ecg693,ecg694,ecg695,ecg696,ecg697,ecg698,ecg699,ecg700,ecg701,ecg702,ecg703,ecg704,ecg705,ecg706,ecg707,ecg708,ecg709,ecg710,ecg711,ecg712,ecg713,ecg714,ecg715,ecg716,ecg717,ecg718,ecg719,ecg720,ecg721,ecg722,ecg723,ecg724,ecg725,ecg726,ecg727,ecg728,ecg729,ecg730,ecg731,ecg732,ecg733,ecg734,ecg735,ecg736,ecg737,ecg738,ecg739,ecg740,ecg741,ecg742,ecg743,ecg744,ecg745,ecg746,ecg747,ecg748,ecg749,ecg750,ecg751,ecg752,ecg753,ecg754,ecg755,ecg756,ecg757,ecg758,ecg759,ecg760,ecg761,ecg762,ecg763,ecg764,ecg765,ecg766,ecg767,ecg768,ecg769,ecg770,ecg771,ecg772,ecg773,ecg774,ecg775,ecg776,ecg777,ecg778,ecg779,ecg780,ecg781,ecg782,ecg783,ecg784,ecg785,ecg786,ecg787,ecg788,ecg789,ecg790,ecg791,ecg792,ecg793,ecg794,ecg795,ecg796,ecg797,ecg798,ecg799,clk,nReset);

endmodule

